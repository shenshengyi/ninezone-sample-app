{"bisBaseClass":"SpatialViewDefinition","viewDefinitionProps":{"classFullName":"BisCore:SpatialViewDefinition","id":"0x70","jsonProperties":{"viewDetails":{"gridOrient":4,"gridPerRef":100,"gridSpaceX":0.1}},"code":{"spec":"0x1c","scope":"0x17","value":"3D Metric Design Model Views - View 1"},"model":"0x17","categorySelectorId":"0x73","displayStyleId":"0x72","isPrivate":false,"description":"","cameraOn":true,"origin":[-70.50636921892303,3.751602553773231,-15.462480803459167],"extents":[107.56996447912394,49.993834494309134,124.11134373851564],"angles":{"pitch":-42.38875364730697,"roll":-55.480840334036685,"yaw":24.87562520991037},"camera":{"lens":46.692503527388425,"focusDist":124.61034373851388,"eye":[-110.70845094680311,-104.99493625015656,59.394984406093556]},"modelSelectorId":"0x71"},"categorySelectorProps":{"classFullName":"BisCore:CategorySelector","id":"0x73","code":{"spec":"0x8","scope":"0x17","value":"3D Metric Design Model Views - View 1"},"model":"0x17","categories":["0x18","0x4f","0x51","0x53","0x55","0x57","0x59","0x5b","0x5d","0x5f","0x61","0x63","0x65","0x67","0x69","0x6b"]},"displayStyleProps":{"classFullName":"BisCore:DisplayStyle3d","id":"0x72","jsonProperties":{"styles":{"hline":{"visible":{"ovrColor":true,"color":0,"pattern":0,"width":1},"hidden":{"ovrColor":true,"color":0,"pattern":3435973836,"width":1},"transThreshold":0.3},"sceneLights":{"ambient":{"intensity":20,"type":2},"sun":{"intensity":99415.46481844832,"type":1},"sunDir":[-6.123233995736766e-17,-3.749399456654644e-33,-1],"portrait":{"intensity":100,"intensity2":100,"type":4},"fstop":0.8570573925971985},"viewflags":{"grid":true,"noSolarLight":true,"noSourceLights":true,"renderMode":6,"visEdges":true},"environment":{"ground":{"aboveColor":32768,"belowColor":1262987,"display":false,"elevation":-0.01},"sky":{"display":false,"groundColor":8228728,"groundExponent":4,"image":{"texture":"0","type":0},"nadirColor":3880,"skyColor":16764303,"skyExponent":4,"zenithColor":16741686}}}},"code":{"spec":"0xa","scope":"0x17","value":"3D Metric Design Model Views - View 1"},"model":"0x17"},"modelSelectorProps":{"classFullName":"BisCore:ModelSelector","id":"0x71","code":{"spec":"0x11","scope":"0x17","value":"3D Metric Design Model Views - View 1"},"model":"0x17","models":["0x40"]}}