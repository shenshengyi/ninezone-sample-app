{"viewDefinitionProps":{"classFullName":"BisCore:SpatialViewDefinition","id":"0x79","jsonProperties":{"viewDetails":{"gridOrient":4,"gridPerRef":100,"gridSpaceX":0.1}},"code":{"spec":"0x1c","scope":"0x17","value":"3D Metric Design Model Views - View 1"},"model":"0x17","categorySelectorId":"0x7c","displayStyleId":"0x7b","isPrivate":false,"description":"","cameraOn":true,"origin":[0.5300491047764453,6.499840034507428,-0.5479192489422662],"extents":[13.271094975461551,5.779961135444573,15.681507674627284],"angles":{"pitch":-42.38875364730822,"roll":-55.48084033403709,"yaw":24.875625209910105},"camera":{"lens":45.87079213591108,"focusDist":15.681507674627259,"eye":[-5.034715583584294,-7.462500355256719,8.849426842976326]},"modelSelectorId":"0x7a"},"categorySelectorProps":{"classFullName":"BisCore:CategorySelector","id":"0x7c","code":{"spec":"0x8","scope":"0x17","value":"3D Metric Design Model Views - View 1"},"model":"0x17","categories":["0x18","0x54","0x56","0x58","0x5a","0x5c","0x5e","0x60","0x62","0x64","0x66","0x68","0x6a","0x6c","0x6e","0x70","0x72","0x74"]},"displayStyleProps":{"classFullName":"BisCore:DisplayStyle3d","id":"0x7b","jsonProperties":{"styles":{"hline":{"visible":{"ovrColor":true,"color":0,"pattern":0,"width":1},"hidden":{"ovrColor":true,"color":0,"pattern":3435973836,"width":1},"transThreshold":0.3},"sceneLights":{"ambient":{"intensity":20,"type":2},"sun":{"intensity":99415.46481844832,"type":1},"sunDir":[-6.123233995736766e-17,-3.749399456654644e-33,-1],"portrait":{"intensity":100,"intensity2":100,"type":4},"fstop":2.9997010231018066},"viewflags":{"grid":true,"noSolarLight":true,"noSourceLights":true,"renderMode":6,"visEdges":true},"environment":{"ground":{"aboveColor":32768,"belowColor":1262987,"display":false,"elevation":-0.01},"sky":{"display":false,"groundColor":8228728,"groundExponent":4,"image":{"texture":"0","type":0},"nadirColor":3880,"skyColor":16764303,"skyExponent":4,"zenithColor":16741686}}}},"code":{"spec":"0xa","scope":"0x17","value":"3D Metric Design Model Views - View 1"},"model":"0x17"},"modelSelectorProps":{"classFullName":"BisCore:ModelSelector","id":"0x7a","code":{"spec":"0x11","scope":"0x17","value":"3D Metric Design Model Views - View 1"},"model":"0x17","models":["0x40"]},"bisBaseClass":"SpatialViewDefinition"}